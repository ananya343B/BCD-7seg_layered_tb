interface intf();
  logic [3:0] s;
  logic [6:0] t;
 
endinterface
